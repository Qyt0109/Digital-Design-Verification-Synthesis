
   reg [8:0] <name> [2047:0]; // 2D 2k * 9
				
				
   wire [2:0] <name>;
				
				
   tri1 [7:0] <name>;
					
					
   // Stores last value when 3-stated
   trireg [1:0] <name> = 2'b00;
						
						