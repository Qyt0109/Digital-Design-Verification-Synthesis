// Convert to a Signed value
$signed(<signal>);
				
				
// Convert to an Unsigned value
$unsigned(<signal>);