// Pause simulation
$stop;
				
// Quit simulation
$finish;