// Assign a value to a signal
assign <reg> = <value>;
			
// Deassign a signal			
deassign <reg>;
			
// Force a signal			
force <wire_or_reg> = <value>;
			
// Release a forced signal
release <wire_or_reg>;

