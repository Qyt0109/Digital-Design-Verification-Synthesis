
/* Multiple lines comment
   Comment here
   Comment here
   Comment here */

// Single line comment
