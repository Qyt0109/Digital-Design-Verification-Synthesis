
#<delay_value>; // Finite delay
			
			
@(<signal>); // Wait for any signal transition
			
			
@(negedge <signal>); // Wait for negative signal transition
			
			
@(posedge <signal>); // Wait for negative signal transition
			
			
wait (<signal>==<value>); // Wait for signal condition
			
		