
<reg> = $random(<seed>);
			
			